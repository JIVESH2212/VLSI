module Decoder_method1(f,x);
	input [3:0] x;
	output reg [15:0] f;
	
	always @(*)
	begin
		if(x == 4'b0000)
			f=16'b0000_0000_0000_0001;
		else if(x == 4'b0001)
			f=16'b0000_0000_0000_0010;
		else if(x == 4'b0010)
			f=16'b0000_0000_0000_0100;
		else if(x == 4'b0011)
			f=16'b0000_0000_0000_1000;
		else if(x == 4'b0100)
			f=16'b0000_0000_0001_0000;
		else if(x == 4'b0101)
			f=16'b0000_0000_0010_0000;
		else if(x == 4'b0110)
			f=16'b0000_0000_0100_0000;
		else if(x == 4'b0111)
			f=16'b0000_0000_1000_0000;
		else if(x == 4'b1000)
			f=16'b0000_0001_0000_0000;
		else if(x == 4'b1001)
			f=16'b0000_0010_0000_0000;
		else if(x == 4'b1010)
			f=16'b0000_0100_0000_0000;
		else if(x == 4'b1011)
			f=16'b0000_1000_0000_0000;
		else if(x == 4'b1100)
			f=16'b0001_0000_0000_0000;
		else if(x == 4'b1101)
			f=16'b0010_0000_0000_0000;
		else if(x == 4'b1110)
			f=16'b0100_0000_0000_0000;
		else if(x == 4'b1111)
			f=16'b1000_0000_0000_0000;
		else //default
			f=16'b0000_0000_0000_0000;
		
	
	end 
	
endmodule
///////////////////////////////////////////////////////
module Decoder_method2(f,x);
	input [3:0] x;
	output reg [15:0] f;
	
	always @(*)
	begin
		case(x)
		4'b0000:
			f=16'b0000_0000_0000_0001;
		4'b0001:
			f=16'b0000_0000_0000_0010;
		4'b0010:
			f=16'b0000_0000_0000_0100;
		4'b0011:
			f=16'b0000_0000_0000_1000;
		4'b0100:
			f=16'b0000_0000_0001_0000;
		4'b0101:
			f=16'b0000_0000_0010_0000;
		4'b0110:
			f=16'b0000_0000_0100_0000;
		4'b0111:
			f=16'b0000_0000_1000_0000;
		4'b1000:
			f=16'b0000_0001_0000_0000;
		4'b1001:
			f=16'b0000_0010_0000_0000;
		4'b1010:
			f=16'b0000_0100_0000_0000;
		4'b1011:
			f=16'b0000_1000_0000_0000;
		4'b1100:
			f=16'b0001_0000_0000_0000;
		4'b1101:
			f=16'b0010_0000_0000_0000;
		4'b1110:
			f=16'b0100_0000_0000_0000;
		4'b1111:
			f=16'b1000_0000_0000_0000;
		default:
			f=16'b0000_0000_0000_0000;
		
		endcase

	end 
	
endmodule

///////////////////////////////////////////////////////
module Decoder_method3(f,x);
	input [3:0] x;
	output wire [15:0] f;
	
	assign f[0] = (~x[3])&(~x[2])&(~x[1])&(~x[0]);
	assign f[1] = (~x[3])&(~x[2])&(~x[1])&(x[0]);
	assign f[2] = (~x[3])&(~x[2])&(x[1])&(~x[0]);
	assign f[3] = (~x[3])&(~x[2])&(x[1])&(x[0]);

	assign f[4] = (~x[3])&(x[2])&(~x[1])&(~x[0]);
	assign f[5] = (~x[3])&(x[2])&(~x[1])&(x[0]);
	assign f[6] = (~x[3])&(x[2])&(x[1])&(~x[0]);
	assign f[7] = (~x[3])&(x[2])&(x[1])&(x[0]);

	assign f[8] = (x[3])&(~x[2])&(~x[1])&(~x[0]);
	assign f[9] = (x[3])&(~x[2])&(~x[1])&(x[0]);
	assign f[10] = (x[3])&(~x[2])&(x[1])&(~x[0]);
	assign f[11] = (x[3])&(~x[2])&(x[1])&(x[0]);

	assign f[12] = (x[3])&(x[2])&(~x[1])&(~x[0]);
	assign f[13] = (x[3])&(x[2])&(~x[1])&(x[0]);
	assign f[14] = (x[3])&(x[2])&(x[1])&(~x[0]);
	assign f[15] = (x[3])&(x[2])&(x[1])&(x[0]);
	
endmodule




///////////////////////////////////////////////////////
module Decoder_method4(f,x);
	input [3:0] x;
	output wire [15:0] f;
	
		assign f = 16'b0000_0000_0000_0001<<x;
	
endmodule